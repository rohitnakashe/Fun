module top_module( 
    input a, 
    input b, 
    output out );

  assign out = a && b; // bitwise-AND (&),  logical-AND (&&) operator

endmodule
