module top_module ( input a, input b, output out );

    mod_a inst1(a , b ,out);
endmodule
